import alu::*;