import ram16::*;

package ram512 (
    input [511:0]in;
    input [8:0]addr;
    input load;
    input clk
    output [511:0]out;
);

wire [15:0]    [511:0]  in0 = in;
wire [31:15]   [511:0]  in1 = in;
wire [47:31]   [511:0]  in2 = in;
wire [63:47]   [511:0]  in3 = in;
wire [79:63]   [511:0]  in4 = in;
wire [95:79]   [511:0]  in5 = in;
wire [111:95]  [511:0]  in6 = in;
wire [127:111] [511:0]  in7 = in;
wire [143:127] [511:0]  in8 = in;
wire [159:143] [511:0]  in9 = in;
wire [179:159] [511:0]  in10 = in;
wire [191:179] [511:0]  in11 = in;
wire [207:191] [511:0]  in12 = in;
wire [223:207] [511:0]  in13 = in;
wire [239:223] [511:0]  in14 = in;
wire [255:239] [511:0]  in15 = in;
wire [271:255] [511:0]  in16 = in;
wire [287:271] [511:0]  in17 = in;
wire [303:287] [511:0]  in18 = in;
wire [319:303] [511:0]  in19 = in;
wire [335:319] [511:0]  in20 = in;
wire [351:335] [511:0]  in21 = in;
wire [367:351] [511:0]  in22 = in;
wire [383:367] [511:0]  in23 = in;
wire [399:383] [511:0]  in24 = in;
wire [415:399] [511:0]  in25 = in;
wire [431:415] [511:0]  in26 = in;
wire [447:431] [511:0]  in27 = in;
wire [463:447] [511:0]  in28 = in;
wire [479:463] [511:0]  in29 = in;
wire [495:479] [511:0]  in30 = in;
wire [511:495] [511:0]  in31 = in;

wire [8:0] [5:0] addr0 = in;
wire [0:8] [5:0] addr1 = in;

wire [15:0]out0;
wire [15:0]out1;
wire [15:0]out2;
wire [15:0]out3;
wire [15:0]out4;
wire [15:0]out5;
wire [15:0]out6;
wire [15:0]out7;
wire [15:0]out8;
wire [15:0]out9;
wire [15:0]out10;
wire [15:0]out11;
wire [15:0]out12;
wire [15:0]out13;
wire [15:0]out14;
wire [15:0]out15;
wire [15:0]out16;
wire [15:0]out17;
wire [15:0]out18;
wire [15:0]out19;
wire [15:0]out20;
wire [15:0]out21;
wire [15:0]out22;
wire [15:0]out23;
wire [15:0]out24;
wire [15:0]out25;
wire [15:0]out26;
wire [15:0]out27;
wire [15:0]out28;
wire [15:0]out29;
wire [15:0]out30;
wire [15:0]out31;

ram16   clstr0(in0, addr0, load, clk, out0);
ram16   clstr1(in1, addr0, load, clk, out1);
ram16   clstr2(in2, addr0, load, clk, out2);
ram16   clstr3(in3, addr0, load, clk, out3);
ram16   clstr4(in4, addr0, load, clk, out4);
ram16   clstr5(in5, addr0, load, clk, out5);
ram16   clstr6(in6, addr0, load, clk, out6);
ram16   clstr7(in7, addr0, load, clk, out7);
ram16   clstr8(in8, addr0, load, clk, out8);
ram16   clstr9(in9, addr0, load, clk, out9);
ram16 clstr10(in10, addr0, load, clk, out10);
ram16 clstr11(in11, addr0, load, clk, out11);
ram16 clstr12(in12, addr0, load, clk, out12);
ram16 clstr13(in13, addr0, load, clk, out13);
ram16 clstr14(in14, addr0, load, clk, out14);
ram16 clstr15(in15, addr0, load, clk, out15);
ram16 clstr16(in16, addr1, load, clk, out16);
ram16 clstr17(in17, addr1, load, clk, out17);
ram16 clstr18(in18, addr1, load, clk, out18);
ram16 clstr19(in19, addr1, load, clk, out19);
ram16 clstr20(in20, addr1, load, clk, out20);
ram16 clstr21(in21, addr1, load, clk, out21);
ram16 clstr22(in22, addr1, load, clk, out22);
ram16 clstr23(in23, addr1, load, clk, out23);
ram16 clstr24(in24, addr1, load, clk, out24);
ram16 clstr25(in25, addr1, load, clk, out25);
ram16 clstr26(in26, addr1, load, clk, out26);
ram16 clstr27(in27, addr1, load, clk, out27);
ram16 clstr28(in28, addr1, load, clk, out28);
ram16 clstr29(in29, addr1, load, clk, out29);
ram16 clstr30(in30, addr1, load, clk, out30);
ram16 clstr31(in31, addr1, load, clk, out31);

wire [15:0]    [511:0]  out0 = out;
wire [31:15]   [511:0]  out1 = out;
wire [47:31]   [511:0]  out2 = out;
wire [63:47]   [511:0]  out3 = out;
wire [79:63]   [511:0]  out4 = out;
wire [95:79]   [511:0]  out5 = out;
wire [111:95]  [511:0]  out6 = out;
wire [127:111] [511:0]  out7 = out;
wire [143:127] [511:0]  out8 = out;
wire [159:143] [511:0]  out9 = out;
wire [179:159] [511:0]  out10 = out;
wire [191:179] [511:0]  out11 = out;
wire [207:191] [511:0]  out12 = out;
wire [223:207] [511:0]  out13 = out;
wire [239:223] [511:0]  out14 = out;
wire [255:239] [511:0]  out15 = out;
wire [271:255] [511:0]  out16 = out;
wire [287:271] [511:0]  out17 = out;
wire [303:287] [511:0]  out18 = out;
wire [319:303] [511:0]  out19 = out;
wire [335:319] [511:0]  out20 = out;
wire [351:335] [511:0]  out21 = out;
wire [367:351] [511:0]  out22 = out;
wire [383:367] [511:0]  out23 = out;
wire [399:383] [511:0]  out24 = out;
wire [415:399] [511:0]  out25 = out;
wire [431:415] [511:0]  out26 = out;
wire [447:431] [511:0]  out27 = out;
wire [463:447] [511:0]  out28 = out;
wire [479:463] [511:0]  out29 = out;
wire [495:479] [511:0]  out30 = out;
wire [511:495] [511:0]  out31 = out;


endpackage