module not16(y16, a16);
    input [15:0] a16;
    output [15:0] y16;

    not(y16[0], a16[0]);
    not(y16[1], a16[1]);
    not(y16[2], a16[2]);
    not(y16[3], a16[3]);
    not(y16[4], a16[4]);
    not(y16[5], a16[5]);
    not(y16[6], a16[6]);
    not(y16[7], a16[7]);
    not(y16[8], a16[8]);
    not(y16[9], a16[9]);
    not(y16[10], a16[10]);
    not(y16[11], a16[11]);
    not(y16[12], a16[12]);
    not(y16[13], a16[13]);
    not(y16[14], a16[14]);
    not(y16[15], a16[15]);
endmodule