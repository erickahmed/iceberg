'`include "gates/"

import name::scope;